module instruction_memory(input wire [31:0] pc,
                          output reg [31:0] instr);

    /*
    L7: lw x6, -4(x9)        I   111111111100 01001 010 00110 0000011
        sw x6, 8(x9)         S   0000000 00110 01001 010 01000 0100011
        or x4, x5, x6        R   0000000 00110 00101 110 00100 0110011
        addi x4, x4, 2       I   000000000010 00100 000 00100 0010011
        and x4, x4, x6       R   0000000 00110 00100 111 00100 0110011
        beq x4, x4, L7       B   1111111 00100 00100 000 01101 1100011

    L8: addi x1, x1, 2       I   000000000010 00001 000 00001 0010011
        and x2, x9, x4       R   0000000 00100 01001 111 00010 0110011
        or x9, x4, x5        R   0000000 00101 00100 110 01001 0110011
        beq x1, x1, L7       B   1111111 00001 00001 000 10101 1100011

            32'h0000: instr = 32'b00000000001000001000000010010011;
            32'h0004: instr = 32'b00000000010001001111000100110011;
            32'h0008: instr = 32'b00000000010100100110010010110011;
            32'h000c: instr = 32'b11111110000100001000101011100011;

    L9: addi x8, x4, 4       I   000000000100 00100 000 01000 0010011
        and x2, x8, x9       R   0000000 01001 01000 111 00010 0110011
        or x3, x4, x8        R   0000000 01000 00100 110 00011 0110011
        and x1, x8, x1       R   0000000 00001 01000 111 00001 0110011
    */

    always @* begin
        case(pc)
            32'h0000: instr = 32'b00000000010000100000010000010011;
            32'h0004: instr = 32'b00000000100101000111000100110011;
            32'h0008: instr = 32'b00000000100000100110000110110011;
            32'h000c: instr = 32'b00000000000101000111000010110011;

            default:  instr = 32'b0;
        endcase
    end
    
endmodule